module regfile(
	input sourceReg1_i,
	input sourceReg2_i,
	input destReg_i,
	input regwrite_i,
	input clk
);